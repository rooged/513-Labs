module Au_32b_tb();

reg[31:0] a,b,s;
reg ALUop;

//wire [31:0] s;

Au_32b ca(.a(a),.b(b),.ALUop(ALUop),.clk(clk),.rst_n(rst_n),.s(s),.hi(hi),.lo(lo),.zero(zero));

initial begin
    #100 a=32'b00000000000000000000000000000001; b=32'b00000000000000000000000000000010; ALUop=2'b00; //sum should be 0011
    #100 a=32'b00000000000000000000000000000010; b=32'b00000000000000000000000000000001; ALUop=2'b01; //sum should be 0001
    #100 a=32'b00000000000000000000000000000011; b=32'b00000000000000000000000000000001; ALUop=2'b00; //sum should be 0100
    #100 a=32'b00000000000000000000000000001000; b=32'b00000000000000000000000000000011; ALUop=2'b01; //sum should be 0101
    #100 a=32'b00000000000000000000000000001000; b=32'b00000000000000000000000000000011; ALUop=2'b00; //sum should be 1011
    #100 a=32'b00000000000000000000000000001010; b=32'b00000000000000000000000000001010; ALUop=2'b01; //sum should be 0000
    #100 a=32'b00000000000000000000000000001010; b=32'b00000000000000000000000000001010; ALUop=2'b00; //sum should be (01)0100
    #100 a=32'b00000000000000000000000000001001; b=32'b00000000000000000000000000000011; ALUop=2'b01; //sum should be 0110
    #100 a=32'b00000000000000000000000000001111; b=32'b00000000000000000000000000000001; ALUop=2'b01; //sum should be 1110
    #100 a=32'b11111111111111111111111111111111; b=32'b00000000000000000000000000000001; ALUop=2'b01;
    #100 a=32'b11111111111111111111111111111111; b=32'b00000000000000000000000000000001; ALUop=2'b00;
    #100 a=32'b11111111111111111111111111111111; b=32'b00000000000000000000000000000011; ALUop=2'b01;
    //#10 $finish;
end
endmodule